module Accelerator(
    input clk, rst, 
    input wStart, lp,
    input [4:0] v,
    input [1:0] u,

    output wrReq, rdReq, wDone
    output [20:0] wrData,
);

    WrapperController()

endmodule